module immediate_selector(
    
)
endmodule;
