module _sll_impl ( // barrel shifter
    input logic [31:0] a,
    input logic [31:0] b,
    output logic [31:0] aer
); 
    always_comb begin
    end

endmodule;