module _slt_impl ( // barrel shifter
    input logic [31:0] a,
    input logic [31:0] b,
    output logic [31:0] aer
); 
    


endmodule;