module sign_extender ( // depreciated/reference
    input logic [24:0] imm_val, // non-extended input
    input logic [2:0] imm_type, // bit source
    output logic [31:0] ext_imm // extended output
)

    always_comb begin
        case (imm_type)
            3'b001: begin // i-type instructions
                as_imm = {{20{imm_val[24]}}, imm_val[24:13]};
            end
            3'b010: begin // s-type instructions
                as_imm = {{20{imm_val[24]}}, imm_val[24:18], imm_val[4:0]}
            end
            3'b011: begin // b-type instructions
                as_imm = {{20{imm_val[24]}}, imm_val[0], imm_val[23:18], imm_val[4:1], 1'b0}
            end
            3'b100: begin // j-type instructions
                as_imm = {{12{imm_val[24]}}, imm_val[12:5], imm_val[13], imm_val[23:14], 1'b0}
            end
            3'b101: begin // u-type instruction (load upper immediate (lui))
                as_imm = {imm_val[24:5], 12{1'b0}};
            end
            default: begin // no immediate
                as_imm = {32{1'b0}};
            end
        endcase
    end

endmodule;